-- Testbench automatically generated online
-- at https://vhdl.lapinoo.net
-- Generation date : 14.6.2023 15:10:21 UTC

library ieee;
use ieee.std_logic_1164.all;
use IEEE.NUMERIC_STD.ALL;
use work.types_pkg.all;

entity teletext_generator_tb is
end teletext_generator_tb;

architecture tb of teletext_generator_tb is

    component teletext_generator
        port (CLK_IN              : in    std_logic;
            RESET_N             : in    std_logic;
            LINE_IN             : in    TELETEXT_LINE;
            PAGE_CONTROL_BITS   : in    CONTROL_BITS;
            PAGE_NUMBER         : in    unsigned (7 downto 0);
            MAGAZINE_NUMBER     : in    unsigned (2 downto 0);
            
            LINE_INDEX          : out   unsigned (4 downto 0);
            
            DATA_OUT            : out   std_logic;
            SYNC_OUT            : out   std_logic
        );
    end component;

    signal CLK_IN   : std_logic;
    signal RESET_N  : std_logic;
    
    signal DATA_OUT : std_logic;
    signal SYNC_OUT : std_logic;
    
    signal LINE_INDEX   : unsigned(4 downto 0);

    constant PAGE_CONTROL_BITS : CONTROL_BITS := (
        ERASE_PAGE => '0',
        NEWSFLASH => '0',
        SUBTITLE => '0',
        SUPPRESS_HEADER => '0',
        UPDATE_INDICATOR => '0',
        INTERRUPTED_SEQUENCE => '0',
        INHIBIT_DISPLAY => '0',
        MAGAZINE_SERIAL => '0',
        NATIONAL_OPTION_CHARACTER_SUBSET => "000"
    );
    constant PAGE_NUMBER : unsigned (7 downto 0) := "00010001";
    
    constant EMPTY_LINE : TELETEXT_LINE := (others => "0100000");

    constant TbPeriod : time := (1000 ns) / 7;
    signal TbClock : std_logic := '0';
    signal TbSimEnded : std_logic := '0';

    signal packet : std_logic_vector (359 downto 0);
    
    signal packet_num: unsigned(4 downto 0);
    signal first_triplet_hamming: std_logic_vector(23 downto 0);
    signal first_hamming_parity: std_logic_vector(5 downto 0);
    signal first_triplet: std_logic_vector(17 downto 0);
    
    signal first_triplet_decoded: TRIPLET;

begin

    dut : teletext_generator
    port map (CLK_IN            => CLK_IN,
              RESET_N           => RESET_N,
              
              LINE_IN           => EMPTY_LINE,
              LINE_INDEX        => LINE_INDEX,
              
              MAGAZINE_NUMBER   => "001",
              
              PAGE_CONTROL_BITS => PAGE_CONTROL_BITS,
              PAGE_NUMBER       => PAGE_NUMBER,
              DATA_OUT          => DATA_OUT,
              SYNC_OUT          => SYNC_OUT);

    -- Clock generation
    TbClock <= not TbClock after TbPeriod/2 when TbSimEnded /= '1' else '0';

    -- EDIT: Check that CLK_IN is really your main clock signal
    CLK_IN <= TbClock;
    
    packet_num <= unsigned(packet(320 downto 320) & packet(322) & packet(324) & packet(326) & packet(328));
    
    first_triplet_hamming <= reverse_any_vector(packet(311 downto 288));
    
    first_triplet <= first_triplet_hamming(22 downto 16) & first_triplet_hamming(14 downto 8) & first_triplet_hamming(6 downto 4) & first_triplet_hamming(2);
    
    first_triplet_decoded.ADDRESS <= unsigned(first_triplet(5 downto 0));
    first_triplet_decoded.MODE <= unsigned(first_triplet(10 downto 6));
    first_triplet_decoded.DATA <= unsigned(first_triplet(17 downto 11));

    first_hamming_parity(0) <= xor (first_triplet_hamming(0 downto 0) & first_triplet_hamming(2) & first_triplet_hamming(4) & first_triplet_hamming(6)
        & first_triplet_hamming(8) & first_triplet_hamming(10) & first_triplet_hamming(12) & first_triplet_hamming(14) 
        & first_triplet_hamming(16) & first_triplet_hamming(18) & first_triplet_hamming(20) & first_triplet_hamming(22));
        
    first_hamming_parity(1) <= xor (first_triplet_hamming(2 downto 1) & first_triplet_hamming(6 downto 5) & first_triplet_hamming(10 downto 9) & first_triplet_hamming(14 downto 13) & first_triplet_hamming(18 downto 17) & first_triplet_hamming(22 downto 21));

    first_hamming_parity(2) <= xor (first_triplet_hamming(6 downto 3) & first_triplet_hamming(14 downto 11) & first_triplet_hamming(22 downto 19));
    
    first_hamming_parity(3) <= xor first_triplet_hamming(14 downto 7);
    
    first_hamming_parity(4) <= xor first_triplet_hamming(22 downto 15);
    
    first_hamming_parity(5) <= xor first_triplet_hamming;

    stimuli : process
    begin
        -- EDIT Adapt initialization as needed

        -- Reset generation
        -- EDIT: Check that RESET_N is really your reset signal
        RESET_N <= '0';
        wait for 100 ns;
        RESET_N <= '1';
        wait for 100 ns;

        
        for k in 0 to 50 loop

            wait until rising_edge(DATA_OUT);
            for i in 359 downto 0 loop
                wait until rising_edge(CLK_IN);
                packet(i) <= DATA_OUT;
                --report std_logic'image(DATA_OUT);
            end loop;
            
            if packet_num = 26 then
                report "Enhancement received!";
                report "First triplet:" & to_hstring(first_triplet);
                report "Address: " & to_string(first_triplet_decoded.ADDRESS) &
                        ", Mode: " & to_string(first_triplet_decoded.MODE) &
                        ", Data: " & to_string(first_triplet_decoded.DATA);
            end if;

            --report std_logic_vector'image(packet);
        end loop;

        -- Stop the clock and hence terminate the simulation
        TbSimEnded <= '1';
        assert false report "end of simulation" severity note;
        
        wait;
    end process;

end tb;